-------------- Forwarding Unit ---------------
LIBRARY ieee;
USE ieee.std_logic_1164.all;
use work.components.all;

ENTITY forwarding_unit is
	port( 
			